interface inter;
  logic a,b;
  logic [3:0]y;
endinterface
