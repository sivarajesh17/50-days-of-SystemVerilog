interface inter;
  logic [7:0]d;
  logic [2:0]q;
endinterface
