interface inter;
  logic a,b,c;
  logic sum,carry;
endinterface
