interface inter;
  logic [3:0]i;
  logic [1:0]s;
  logic y;
endinterface
