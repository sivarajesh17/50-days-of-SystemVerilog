interface inter;
  logic din;
  logic [1:0]sel;
  logic [3:0]y;
endinterface
