interface dff_if;
    logic clk;
    logic reset;
    logic d;
    logic q;
endinterface

