interface inter;
  logic [3:0]a,b;
  logic a_gt_b,a_lt_b,a_eq_b;
endinterface

