interface inter;
  logic a,b;
  logic sum,carry;
endinterface
