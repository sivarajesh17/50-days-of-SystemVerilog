interface inter;
  logic [3:0]a,b;
  logic [3:0]sum;
  logic c;
  logic carry;
endinterface
